library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CSA16 is
end CSA16;

architecture Behavioral of CSA16 is

begin


end Behavioral;

